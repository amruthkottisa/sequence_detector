module 
  

module sd(input clk, input rst, input in, output reg out);
  reg [2:0] ps,ns;
  parameter s0=0, 
  
